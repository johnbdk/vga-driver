module VRAM(DIA_R, DIA_G, DIA_B, ADDRA, CLKA, ENA, SSRA, WEA, DOA_R, DOA_G, DOA_B);
input 	DIA_R, DIA_G, DIA_B, ADDRA, CLKA, ENA, SSRA, WEA;
output 	DOA_R, DOA_G, DOA_B;

/* RED COLOR MEMORY */
RAMB16_S1_S1 #(
      .INIT_A(1'b0),                // Value of output RAM registers on Port A at startup
      .INIT_B(1'b0),                // Value of output RAM registers on Port B at startup
      .SRVAL_A(1'b0),               // Port A output value upon SSR assertion
      .SRVAL_B(1'b0),               // Port B output value upon SSR assertion
      .WRITE_MODE_A("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
      .WRITE_MODE_B("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
      .SIM_COLLISION_CHECK("ALL"),  // "NONE", "WARNING_ONLY", "GENERATE_X_ONLY", "ALL" 

      // Address 0 to 4095
      .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_01(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_03(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_05(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_07(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_09(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0B(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0D(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0F(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      // Address 4096 to 8191
      .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 8192 to 12287
      .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 12288 to 16383
      .INIT_30(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_31(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_32(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_33(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_34(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_35(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_36(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_37(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_38(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_39(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_3A(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_3B(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_3C(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_3D(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_3E(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_3F(256'h4444444444444444444444444444444444444444444444444444444444444444)
) RAMB16_S1_S1_red (
      .DOA(DOA_R),      // Port A 1-bit Data Output
      //.DOB(DOB),      // Port B 1-bit Data Output
      .ADDRA(ADDRA),  // Port A 14-bit Address Input
      //.ADDRB(ADDRB),  // Port B 14-bit Address Input
      .CLKA(CLKA),    // Port A Clock
      //.CLKB(CLKB),    // Port B Clock
      .DIA(DIA_R),        // Port A 1-bit Data Input
      //.DIB(DIB),      // Port B 1-bit Data Input
      .ENA(ENA),      // Port A RAM Enable Input
      //.ENB(ENB),      // Port B RAM Enable Input
      .SSRA(SSRA),    // Port A Synchronous Set/Reset Input
      //.SSRB(SSRB),    // Port B Synchronous Set/Reset Input
      .WEA(WEA)      // Port A Write Enable Input
      //.WEB(WEB)       // Port B Write Enable Input
);

/* GREEN COLOR MEMORY */
RAMB16_S1_S1 #(
      .INIT_A(1'b0),                // Value of output RAM registers on Port A at startup
      .INIT_B(1'b0),                // Value of output RAM registers on Port B at startup
      .SRVAL_A(1'b0),               // Port A output value upon SSR assertion
      .SRVAL_B(1'b0),               // Port B output value upon SSR assertion
      .WRITE_MODE_A("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
      .WRITE_MODE_B("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
      .SIM_COLLISION_CHECK("ALL"),  // "NONE", "WARNING_ONLY", "GENERATE_X_ONLY", "ALL" 

      // Address 0 to 4095
      .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 4096 to 8191
      .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_11(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_13(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_15(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_17(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_19(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1B(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1D(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1F(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      // Address 8192 to 12287
      .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 12288 to 16383
      .INIT_30(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_31(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_32(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_33(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_34(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_35(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_36(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_37(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_38(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_39(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_3A(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_3B(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_3C(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_3D(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_3E(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_3F(256'h2222222222222222222222222222222222222222222222222222222222222222)
) RAMB16_S1_S1_green (
      .DOA(DOA_G),      // Port A 1-bit Data Output
      //.DOB(DOB),      // Port B 1-bit Data Output
      .ADDRA(ADDRA),  // Port A 14-bit Address Input
      //.ADDRB(ADDRB),  // Port B 14-bit Address Input
      .CLKA(CLKA),    // Port A Clock
      //.CLKB(CLKB),    // Port B Clock
      .DIA(DIA_G),      // Port A 1-bit Data Input
      //.DIB(DIB),      // Port B 1-bit Data Input
      .ENA(ENA),      // Port A RAM Enable Input
      //.ENB(ENB),      // Port B RAM Enable Input
      .SSRA(SSRA),    // Port A Synchronous Set/Reset Input
      //.SSRB(SSRB),    // Port B Synchronous Set/Reset Input
      .WEA(WEA)      // Port A Write Enable Input
      //.WEB(WEB)       // Port B Write Enable Input
);

/* BLUE COLOR MEMORY */
RAMB16_S1_S1 #(
      .INIT_A(1'b0),                // Value of output RAM registers on Port A at startup
      .INIT_B(1'b0),                // Value of output RAM registers on Port B at startup
      .SRVAL_A(1'b0),               // Port A output value upon SSR assertion
      .SRVAL_B(1'b0),               // Port B output value upon SSR assertion
      .WRITE_MODE_A("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
      .WRITE_MODE_B("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
      .SIM_COLLISION_CHECK("ALL"),  // "NONE", "WARNING_ONLY", "GENERATE_X_ONLY", "ALL" 

      // Address 0 to 4095
      .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 4096 to 8191
      .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 8192 to 12287
      .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_21(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_23(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_25(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_27(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_29(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2B(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2D(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2F(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      // Address 12288 to 16383
      .INIT_30(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_31(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_32(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_33(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_34(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_35(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_36(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_37(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_38(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_39(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_3A(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_3B(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_3C(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_3D(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_3E(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_3F(256'h1111111111111111111111111111111111111111111111111111111111111111)
) RAMB16_S1_S1_blue (
      .DOA(DOA_B),      // Port A 1-bit Data Output
      //.DOB(DOB),      // Port B 1-bit Data Output
      .ADDRA(ADDRA),  // Port A 14-bit Address Input
      //.ADDRB(ADDRB),  // Port B 14-bit Address Input
      .CLKA(CLKA),    // Port A Clock
      //.CLKB(CLKB),    // Port B Clock
      .DIA(DIA_B),      // Port A 1-bit Data Input
      //.DIB(DIB),      // Port B 1-bit Data Input
      .ENA(ENA),      // Port A RAM Enable Input
      //.ENB(ENB),      // Port B RAM Enable Input
      .SSRA(SSRA),    // Port A Synchronous Set/Reset Input
      //.SSRB(SSRB),    // Port B Synchronous Set/Reset Input
      .WEA(WEA)      // Port A Write Enable Input
      //.WEB(WEB)       // Port B Write Enable Input
);

endmodule