module VRAM(DIA_R, DIA_G, DIA_B, ADDRA, clk, ENA, SSRA, WEA, DOA_R, DOA_G, DOA_B);

input       [13:0] ADDRA;
input 	DIA_R, DIA_G, DIA_B, clk, ENA, SSRA, WEA;
output 	DOA_R, DOA_G, DOA_B;

/*    128x96
	24	red lines
	24	blue lines
	24	green lines
	24	mixed vetical
	since block size is 256 bits we need 12 lines of 256 bits (or 64 hex digits)
	where	32	hex digits represent a line (128bits) 
*/
	
/* RED COLOR MEMORY */
   RAMB16_S1 #(
      .INIT(1'b1),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("NO_CHANGE"), // WRITE_FIRST, NO_CHANGE or READ_FIRST

      // Address 0 to 4095
      .INIT_00(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_01(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_02(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_03(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_04(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_05(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_06(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_07(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_08(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_09(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_0A(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_0B(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),//end of 1/4
      .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 4096 to 8191
      .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),//end of 2/4
      .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 8192 to 12287
      .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),//end of 3/4
      .INIT_24(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_25(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_26(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_27(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_28(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_29(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_2A(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_2B(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_2C(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_2D(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_2E(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_2F(256'h4444444444444444444444444444444444444444444444444444444444444444),//end of 4/4
      // Address 12288 to 16383	, not needed
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) RAMB16_S1_inst_red (
      .DO(DOA_R),      // 1-bit Data Output
      .ADDR(ADDRA),  // 14-bit Address Input
      .CLK(clk),    // Clock
      .DI(DIA_R),      // 1-bit Data Input
      .EN(ENA),      // RAM Enable Input
      .SSR(SSRA),    // Synchronous Set/Reset Input
      .WE(WEA)       // Write Enable Input
   );

/* GREEN COLOR MEMORY */
   RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("NO_CHANGE"), // WRITE_FIRST, NO_CHANGE or READ_FIRST

      // Address 0 to 4095
      .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),//end of 1/4
      .INIT_0C(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_0D(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_0E(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_0F(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      // Address 4096 to 8191
      .INIT_10(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_11(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_12(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_13(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_14(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_15(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_16(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_17(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),//end of 2/4
      .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 8192 to 12287
      .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),//end of 3/4
      .INIT_24(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_25(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_26(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_27(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_28(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_29(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_2A(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_2B(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_2C(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_2D(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_2E(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_2F(256'h2222222222222222222222222222222222222222222222222222222222222222),//end of 4/4
      // Address 12288 to 16383
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) RAMB16_S1_inst_green (
      .DO(DOA_G),      // 1-bit Data Output
      .ADDR(ADDRA),  // 14-bit Address Input
      .CLK(clk),    // Clock
      .DI(DIA_G),      // 1-bit Data Input
      .EN(ENA),      // RAM Enable Input
      .SSR(SSRA),    // Synchronous Set/Reset Input
      .WE(WEA)       // Write Enable Input
   );

/* BLUE COLOR MEMORY */
   RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("NO_CHANGE"), // WRITE_FIRST, NO_CHANGE or READ_FIRST

      // Address 0 to 4095
      .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),//end of 1/4
      .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 4096 to 8191
      .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),//end of 2/4
      .INIT_18(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_19(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_1A(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_1B(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_1C(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_1D(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_1E(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_1F(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      // Address 8192 to 12287
      .INIT_20(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_21(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_22(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),
      .INIT_23(256'h00000000000000000000000000000000ffffffffffffffffffffffffffffffff),//end of 3/4
      .INIT_24(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_25(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_26(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_27(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_28(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_29(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_2A(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_2B(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_2C(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_2D(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_2E(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_2F(256'h1111111111111111111111111111111111111111111111111111111111111111),//end of 4/4
      // Address 12288 to 16383
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) RAMB16_S1_inst_blue (
      .DO(DOA_B),      // 1-bit Data Output
      .ADDR(ADDRA),  // 14-bit Address Input
      .CLK(clk),    // Clock
      .DI(DIA_B),      // 1-bit Data Input
      .EN(ENA),      // RAM Enable Input
      .SSR(SSRA),    // Synchronous Set/Reset Input
      .WE(WEA)      // Write Enable Input
   );

endmodule